library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 13;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : std_logic_vector(3 downto 0) := "1001";
  constant RET  : std_logic_vector(3 downto 0) := "1010";
  constant ANDOP: std_logic_vector(3 downto 0) := "1011";
  constant ADDI : std_logic_vector(3 downto 0) := "1100";
  constant SUBI : std_logic_vector(3 downto 0) := "1101";
  constant ANDI : std_logic_vector(3 downto 0) := "1110";

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
      -- Inicializa os endereços:
tmp(0) := LDI&"00"&'0'&x"00";
tmp(1) := STA&"00"&'1'&x"20";
tmp(2) := STA&"00"&'1'&x"21";
tmp(3) := STA&"00"&'1'&x"22";
tmp(4) := STA&"00"&'1'&x"23";
tmp(5) := STA&"00"&'1'&x"24";
tmp(6) := STA&"00"&'1'&x"25";
tmp(7) := STA&"00"&'1'&x"00";
tmp(8) := STA&"00"&'1'&x"01";
tmp(9) := STA&"00"&'1'&x"02";
tmp(10) := STA&"00"&'0'&x"00";
tmp(11) := STA&"00"&'0'&x"01";
tmp(12) := STA&"00"&'0'&x"02";
tmp(13) := STA&"00"&'0'&x"03";
tmp(14) := STA&"00"&'0'&x"04";
tmp(15) := STA&"00"&'0'&x"05";
tmp(16) := STA&"00"&'0'&x"06";
tmp(17) := STA&"00"&'1'&x"ff";
tmp(18) := STA&"00"&'1'&x"fe";
tmp(19) := LDI&"00"&'0'&x"01";
tmp(20) := STA&"00"&'0'&x"0e";
tmp(21) := LDI&"00"&'0'&x"0a";
tmp(22) := STA&"00"&'0'&x"0f";
tmp(23) := LDI&"00"&'0'&x"00";
tmp(24) := STA&"00"&'0'&x"10";
tmp(25) := LDI&"00"&'0'&x"06";
tmp(26) := STA&"00"&'0'&x"11";
tmp(27) := LDI&"00"&'0'&x"09";
tmp(28) := STA&"00"&'0'&x"08";
tmp(29) := STA&"00"&'0'&x"0a";
tmp(30) := LDI&"00"&'0'&x"05";
tmp(31) := STA&"00"&'0'&x"09";
tmp(32) := STA&"00"&'0'&x"0b";
tmp(33) := LDI&"00"&'0'&x"03";
tmp(34) := STA&"00"&'0'&x"0c";
tmp(35) := LDI&"00"&'0'&x"02";
tmp(36) := STA&"00"&'0'&x"0d";
tmp(38) := LDI&"00"&'0'&x"0a";
tmp(39) := STA&"00"&'0'&x"12";
tmp(40) := STA&"00"&'0'&x"13";
tmp(41) := STA&"00"&'0'&x"14";
tmp(42) := STA&"00"&'0'&x"15";
tmp(43) := STA&"00"&'0'&x"16";
tmp(44) := STA&"00"&'0'&x"17";
tmp(46) := JSR&"00"&'0'&x"44";
tmp(47) := LDA&"00"&'1'&x"60";
tmp(48) := ANDOP&"00"&'0'&x"0e";
tmp(49) := CEQ&"00"&'0'&x"06";
tmp(50) := JEQ&"00"&'0'&x"34";
tmp(51) := JSR&"00"&'0'&x"fa";
tmp(53) := LDA&"00"&'1'&x"61";
tmp(54) := ANDOP&"00"&'0'&x"0e";
tmp(55) := CEQ&"00"&'0'&x"06";
tmp(56) := JEQ&"00"&'0'&x"3a";
tmp(57) := JSR&"00"&'0'&x"9d";
tmp(59) := JSR&"00"&'1'&x"6d";
tmp(60) := JSR&"00"&'1'&x"3e";
tmp(61) := JSR&"00"&'0'&x"57";
tmp(62) := LDA&"00"&'0'&x"10";
tmp(63) := CEQ&"00"&'0'&x"06";
tmp(64) := JEQ&"00"&'0'&x"42";
tmp(65) := JSR&"00"&'1'&x"9d";
tmp(67) := JMP&"00"&'0'&x"2d";
tmp(69) := LDA&"10"&'0'&x"00";
tmp(70) := STA&"10"&'1'&x"20";
tmp(71) := NOP&"00"&'0'&x"00";
tmp(72) := LDA&"10"&'0'&x"01";
tmp(73) := STA&"10"&'1'&x"21";
tmp(74) := NOP&"00"&'0'&x"00";
tmp(75) := LDA&"10"&'0'&x"02";
tmp(76) := STA&"10"&'1'&x"22";
tmp(77) := NOP&"00"&'0'&x"00";
tmp(78) := LDA&"10"&'0'&x"03";
tmp(79) := STA&"10"&'1'&x"23";
tmp(80) := NOP&"00"&'0'&x"00";
tmp(81) := LDA&"10"&'0'&x"04";
tmp(82) := STA&"10"&'1'&x"24";
tmp(83) := NOP&"00"&'0'&x"00";
tmp(84) := LDA&"10"&'0'&x"05";
tmp(85) := STA&"10"&'1'&x"25";
tmp(86) := RET&"00"&'0'&x"00";
tmp(88) := STA&"00"&'1'&x"ff";
tmp(89) := LDA&"00"&'0'&x"10";
tmp(90) := CEQ&"00"&'0'&x"0e";
tmp(91) := JEQ&"00"&'0'&x"9b";
tmp(92) := LDA&"00"&'0'&x"00";
tmp(93) := SOMA&"00"&'0'&x"0e";
tmp(94) := STA&"00"&'0'&x"00";
tmp(95) := CEQ&"00"&'0'&x"0f";
tmp(96) := JEQ&"00"&'0'&x"63";
tmp(97) := NOP&"00"&'0'&x"00";
tmp(98) := RET&"00"&'0'&x"00";
tmp(100) := LDI&"00"&'0'&x"00";
tmp(101) := STA&"00"&'0'&x"00";
tmp(102) := LDA&"00"&'0'&x"01";
tmp(103) := SOMA&"00"&'0'&x"0e";
tmp(104) := STA&"00"&'0'&x"01";
tmp(105) := CEQ&"00"&'0'&x"11";
tmp(106) := JEQ&"00"&'0'&x"6d";
tmp(107) := NOP&"00"&'0'&x"00";
tmp(108) := RET&"00"&'0'&x"00";
tmp(110) := LDI&"00"&'0'&x"00";
tmp(111) := STA&"00"&'0'&x"01";
tmp(112) := LDA&"00"&'0'&x"02";
tmp(113) := SOMA&"00"&'0'&x"0e";
tmp(114) := STA&"00"&'0'&x"02";
tmp(115) := CEQ&"00"&'0'&x"0f";
tmp(116) := JEQ&"00"&'0'&x"77";
tmp(117) := NOP&"00"&'0'&x"00";
tmp(118) := RET&"00"&'0'&x"00";
tmp(120) := LDI&"00"&'0'&x"00";
tmp(121) := STA&"00"&'0'&x"02";
tmp(122) := LDA&"00"&'0'&x"03";
tmp(123) := SOMA&"00"&'0'&x"0e";
tmp(124) := STA&"00"&'0'&x"03";
tmp(125) := CEQ&"00"&'0'&x"11";
tmp(126) := JEQ&"00"&'0'&x"81";
tmp(127) := NOP&"00"&'0'&x"00";
tmp(128) := RET&"00"&'0'&x"00";
tmp(130) := LDI&"00"&'0'&x"00";
tmp(131) := STA&"00"&'0'&x"03";
tmp(132) := LDA&"00"&'0'&x"04";
tmp(133) := SOMA&"00"&'0'&x"0e";
tmp(134) := STA&"00"&'0'&x"04";
tmp(135) := CEQ&"00"&'0'&x"0f";
tmp(136) := JEQ&"00"&'0'&x"8b";
tmp(137) := NOP&"00"&'0'&x"00";
tmp(138) := RET&"00"&'0'&x"00";
tmp(140) := LDI&"00"&'0'&x"00";
tmp(141) := STA&"00"&'0'&x"04";
tmp(142) := LDA&"00"&'0'&x"05";
tmp(143) := SOMA&"00"&'0'&x"0e";
tmp(144) := STA&"00"&'0'&x"05";
tmp(145) := CEQ&"00"&'0'&x"11";
tmp(146) := JEQ&"00"&'0'&x"95";
tmp(147) := NOP&"00"&'0'&x"00";
tmp(148) := RET&"00"&'0'&x"00";
tmp(150) := LDI&"00"&'0'&x"00";
tmp(151) := STA&"00"&'0'&x"05";
tmp(152) := LDI&"00"&'0'&x"01";
tmp(153) := STA&"00"&'1'&x"02";
tmp(154) := STA&"00"&'0'&x"10";
tmp(156) := RET&"00"&'0'&x"00";
tmp(158) := STA&"00"&'1'&x"fe";
tmp(159) := LDI&"01"&'0'&x"00";
tmp(160) := STA&"01"&'1'&x"20";
tmp(161) := STA&"01"&'1'&x"21";
tmp(162) := STA&"01"&'1'&x"22";
tmp(163) := STA&"01"&'1'&x"23";
tmp(164) := STA&"01"&'1'&x"24";
tmp(165) := STA&"01"&'1'&x"25";
tmp(166) := LDI&"00"&'0'&x"01";
tmp(167) := STA&"00"&'1'&x"01";
tmp(168) := STA&"00"&'1'&x"02";
tmp(170) := LDI&"00"&'0'&x"01";
tmp(171) := STA&"00"&'1'&x"00";
tmp(172) := LDA&"00"&'1'&x"40";
tmp(173) := STA&"00"&'0'&x"00";
tmp(174) := STA&"00"&'1'&x"20";
tmp(175) := LDA&"00"&'1'&x"61";
tmp(176) := ANDOP&"00"&'0'&x"0e";
tmp(177) := CEQ&"00"&'0'&x"06";
tmp(178) := JEQ&"00"&'0'&x"a9";
tmp(179) := LDI&"00"&'0'&x"00";
tmp(180) := STA&"00"&'1'&x"00";
tmp(181) := STA&"00"&'1'&x"fe";
tmp(183) := LDI&"00"&'0'&x"02";
tmp(184) := STA&"00"&'1'&x"00";
tmp(185) := LDA&"00"&'1'&x"40";
tmp(186) := STA&"00"&'0'&x"01";
tmp(187) := STA&"00"&'1'&x"21";
tmp(188) := LDA&"00"&'1'&x"61";
tmp(189) := ANDOP&"00"&'0'&x"0e";
tmp(190) := CEQ&"00"&'0'&x"06";
tmp(191) := JEQ&"00"&'0'&x"b6";
tmp(192) := LDI&"00"&'0'&x"00";
tmp(193) := STA&"00"&'1'&x"00";
tmp(194) := STA&"00"&'1'&x"fe";
tmp(196) := LDI&"00"&'0'&x"04";
tmp(197) := STA&"00"&'1'&x"00";
tmp(198) := LDA&"00"&'1'&x"40";
tmp(199) := STA&"00"&'0'&x"02";
tmp(200) := STA&"00"&'1'&x"22";
tmp(201) := LDA&"00"&'1'&x"61";
tmp(202) := ANDOP&"00"&'0'&x"0e";
tmp(203) := CEQ&"00"&'0'&x"06";
tmp(204) := JEQ&"00"&'0'&x"c3";
tmp(205) := LDI&"00"&'0'&x"00";
tmp(206) := STA&"00"&'1'&x"00";
tmp(207) := STA&"00"&'1'&x"fe";
tmp(209) := LDI&"00"&'0'&x"08";
tmp(210) := STA&"00"&'1'&x"00";
tmp(211) := LDA&"00"&'1'&x"40";
tmp(212) := STA&"00"&'0'&x"03";
tmp(213) := STA&"00"&'1'&x"23";
tmp(214) := LDA&"00"&'1'&x"61";
tmp(215) := ANDOP&"00"&'0'&x"0e";
tmp(216) := CEQ&"00"&'0'&x"06";
tmp(217) := JEQ&"00"&'0'&x"d0";
tmp(218) := LDI&"00"&'0'&x"00";
tmp(219) := STA&"00"&'1'&x"00";
tmp(220) := STA&"00"&'1'&x"fe";
tmp(222) := LDI&"00"&'0'&x"10";
tmp(223) := STA&"00"&'1'&x"00";
tmp(224) := LDA&"00"&'1'&x"40";
tmp(225) := STA&"00"&'0'&x"04";
tmp(226) := STA&"00"&'1'&x"24";
tmp(227) := LDA&"00"&'1'&x"61";
tmp(228) := ANDOP&"00"&'0'&x"0e";
tmp(229) := CEQ&"00"&'0'&x"06";
tmp(230) := JEQ&"00"&'0'&x"dd";
tmp(231) := LDI&"00"&'0'&x"00";
tmp(232) := STA&"00"&'1'&x"00";
tmp(233) := STA&"00"&'1'&x"fe";
tmp(235) := LDI&"00"&'0'&x"20";
tmp(236) := STA&"00"&'1'&x"00";
tmp(237) := LDA&"00"&'1'&x"40";
tmp(238) := STA&"00"&'0'&x"05";
tmp(239) := STA&"00"&'1'&x"25";
tmp(240) := LDA&"00"&'1'&x"61";
tmp(241) := ANDOP&"00"&'0'&x"0e";
tmp(242) := CEQ&"00"&'0'&x"06";
tmp(243) := JEQ&"00"&'0'&x"ea";
tmp(244) := LDI&"00"&'0'&x"00";
tmp(245) := STA&"00"&'1'&x"00";
tmp(246) := STA&"00"&'1'&x"fe";
tmp(247) := STA&"00"&'1'&x"01";
tmp(248) := STA&"00"&'1'&x"02";
tmp(249) := RET&"00"&'0'&x"00";
tmp(251) := STA&"00"&'1'&x"ff";
tmp(252) := LDI&"00"&'0'&x"aa";
tmp(253) := STA&"00"&'1'&x"00";
tmp(254) := LDI&"01"&'0'&x"00";
tmp(255) := STA&"01"&'1'&x"20";
tmp(256) := STA&"01"&'1'&x"21";
tmp(257) := STA&"01"&'1'&x"22";
tmp(258) := STA&"01"&'1'&x"23";
tmp(259) := STA&"01"&'1'&x"24";
tmp(260) := STA&"01"&'1'&x"25";
tmp(262) := LDA&"00"&'1'&x"40";
tmp(263) := STA&"00"&'0'&x"12";
tmp(264) := STA&"00"&'1'&x"20";
tmp(265) := LDA&"00"&'1'&x"60";
tmp(266) := ANDOP&"00"&'0'&x"0e";
tmp(267) := CEQ&"00"&'0'&x"06";
tmp(268) := JEQ&"00"&'1'&x"05";
tmp(269) := STA&"00"&'1'&x"ff";
tmp(271) := LDA&"00"&'1'&x"40";
tmp(272) := STA&"00"&'0'&x"13";
tmp(273) := STA&"00"&'1'&x"21";
tmp(274) := LDA&"00"&'1'&x"60";
tmp(275) := ANDOP&"00"&'0'&x"0e";
tmp(276) := CEQ&"00"&'0'&x"06";
tmp(277) := JEQ&"00"&'1'&x"0e";
tmp(278) := STA&"00"&'1'&x"ff";
tmp(280) := LDA&"00"&'1'&x"40";
tmp(281) := STA&"00"&'0'&x"14";
tmp(282) := STA&"00"&'1'&x"22";
tmp(283) := LDA&"00"&'1'&x"60";
tmp(284) := ANDOP&"00"&'0'&x"0e";
tmp(285) := CEQ&"00"&'0'&x"06";
tmp(286) := JEQ&"00"&'1'&x"17";
tmp(287) := STA&"00"&'1'&x"ff";
tmp(289) := LDA&"00"&'1'&x"40";
tmp(290) := STA&"00"&'0'&x"15";
tmp(291) := STA&"00"&'1'&x"23";
tmp(292) := LDA&"00"&'1'&x"60";
tmp(293) := ANDOP&"00"&'0'&x"0e";
tmp(294) := CEQ&"00"&'0'&x"06";
tmp(295) := JEQ&"00"&'1'&x"20";
tmp(296) := STA&"00"&'1'&x"ff";
tmp(298) := LDA&"00"&'1'&x"40";
tmp(299) := STA&"00"&'0'&x"16";
tmp(300) := STA&"00"&'1'&x"24";
tmp(301) := LDA&"00"&'1'&x"60";
tmp(302) := ANDOP&"00"&'0'&x"0e";
tmp(303) := CEQ&"00"&'0'&x"06";
tmp(304) := JEQ&"00"&'1'&x"29";
tmp(305) := STA&"00"&'1'&x"ff";
tmp(307) := LDA&"00"&'1'&x"40";
tmp(308) := STA&"00"&'0'&x"17";
tmp(309) := STA&"00"&'1'&x"25";
tmp(310) := LDA&"00"&'1'&x"60";
tmp(311) := ANDOP&"00"&'0'&x"0e";
tmp(312) := CEQ&"00"&'0'&x"06";
tmp(313) := JEQ&"00"&'1'&x"32";
tmp(314) := LDI&"00"&'0'&x"00";
tmp(315) := STA&"00"&'1'&x"00";
tmp(316) := STA&"00"&'1'&x"ff";
tmp(317) := RET&"00"&'0'&x"00";
tmp(319) := LDA&"01"&'0'&x"05";
tmp(320) := CEQ&"01"&'0'&x"0d";
tmp(321) := JEQ&"00"&'1'&x"45";
tmp(322) := LDI&"01"&'0'&x"00";
tmp(323) := STA&"01"&'0'&x"10";
tmp(324) := RET&"00"&'0'&x"00";
tmp(326) := LDA&"01"&'0'&x"04";
tmp(327) := CEQ&"01"&'0'&x"0c";
tmp(328) := JEQ&"00"&'1'&x"4c";
tmp(329) := LDI&"01"&'0'&x"00";
tmp(330) := STA&"01"&'0'&x"10";
tmp(331) := RET&"00"&'0'&x"00";
tmp(333) := LDA&"01"&'0'&x"03";
tmp(334) := CEQ&"01"&'0'&x"0b";
tmp(335) := JEQ&"00"&'1'&x"53";
tmp(336) := LDI&"01"&'0'&x"00";
tmp(337) := STA&"01"&'0'&x"10";
tmp(338) := RET&"00"&'0'&x"00";
tmp(340) := LDA&"01"&'0'&x"02";
tmp(341) := CEQ&"01"&'0'&x"0a";
tmp(342) := JEQ&"00"&'1'&x"5a";
tmp(343) := LDI&"01"&'0'&x"00";
tmp(344) := STA&"01"&'0'&x"10";
tmp(345) := RET&"00"&'0'&x"00";
tmp(347) := LDA&"01"&'0'&x"01";
tmp(348) := CEQ&"01"&'0'&x"09";
tmp(349) := JEQ&"00"&'1'&x"61";
tmp(350) := LDI&"01"&'0'&x"00";
tmp(351) := STA&"01"&'0'&x"10";
tmp(352) := RET&"00"&'0'&x"00";
tmp(354) := LDA&"01"&'0'&x"00";
tmp(355) := CEQ&"01"&'0'&x"08";
tmp(356) := JEQ&"00"&'1'&x"68";
tmp(357) := LDI&"01"&'0'&x"00";
tmp(358) := STA&"01"&'0'&x"10";
tmp(359) := RET&"00"&'0'&x"00";
tmp(361) := LDI&"01"&'0'&x"01";
tmp(362) := STA&"01"&'0'&x"10";
tmp(363) := STA&"01"&'1'&x"01";
tmp(364) := RET&"00"&'0'&x"00";
tmp(366) := LDA&"01"&'0'&x"05";
tmp(367) := CEQ&"01"&'0'&x"17";
tmp(368) := JEQ&"00"&'1'&x"72";
tmp(369) := RET&"00"&'0'&x"00";
tmp(371) := LDA&"01"&'0'&x"04";
tmp(372) := CEQ&"01"&'0'&x"16";
tmp(373) := JEQ&"00"&'1'&x"77";
tmp(374) := RET&"00"&'0'&x"00";
tmp(376) := LDA&"01"&'0'&x"03";
tmp(377) := CEQ&"01"&'0'&x"15";
tmp(378) := JEQ&"00"&'1'&x"7c";
tmp(379) := RET&"00"&'0'&x"00";
tmp(381) := LDA&"01"&'0'&x"02";
tmp(382) := CEQ&"01"&'0'&x"14";
tmp(383) := JEQ&"00"&'1'&x"81";
tmp(384) := RET&"00"&'0'&x"00";
tmp(386) := LDA&"01"&'0'&x"01";
tmp(387) := CEQ&"01"&'0'&x"13";
tmp(388) := JEQ&"00"&'1'&x"86";
tmp(389) := RET&"00"&'0'&x"00";
tmp(391) := LDA&"01"&'0'&x"00";
tmp(392) := CEQ&"01"&'0'&x"12";
tmp(393) := JEQ&"00"&'1'&x"8b";
tmp(394) := RET&"00"&'0'&x"00";
tmp(396) := LDI&"00"&'0'&x"00";
tmp(397) := LDI&"10"&'0'&x"aa";
tmp(398) := LDI&"01"&'0'&x"55";
tmp(399) := STA&"00"&'1'&x"00";
tmp(400) := NOP&"00"&'0'&x"00";
tmp(401) := STA&"10"&'1'&x"00";
tmp(402) := NOP&"00"&'0'&x"00";
tmp(403) := STA&"00"&'1'&x"00";
tmp(404) := NOP&"00"&'0'&x"00";
tmp(405) := STA&"01"&'1'&x"00";
tmp(406) := LDA&"00"&'1'&x"64";
tmp(407) := ANDOP&"00"&'0'&x"0e";
tmp(408) := CEQ&"00"&'0'&x"06";
tmp(409) := JEQ&"00"&'1'&x"8b";
tmp(410) := STA&"00"&'1'&x"fc";
tmp(411) := STA&"00"&'1'&x"00";
tmp(412) := RET&"00"&'0'&x"00";
tmp(414) := LDI&"00"&'0'&x"00";
tmp(415) := STA&"00"&'0'&x"00";
tmp(416) := STA&"00"&'0'&x"01";
tmp(417) := STA&"00"&'0'&x"02";
tmp(418) := STA&"00"&'0'&x"03";
tmp(419) := STA&"00"&'0'&x"04";
tmp(420) := STA&"00"&'0'&x"05";
tmp(421) := STA&"00"&'0'&x"10";
tmp(422) := STA&"00"&'1'&x"01";
tmp(423) := STA&"00"&'1'&x"02";
tmp(424) := STA&"00"&'1'&x"00";
tmp(425) := RET&"00"&'0'&x"00";





        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;