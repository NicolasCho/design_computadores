library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 13;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : std_logic_vector(3 downto 0) := "1001";
  constant RET  : std_logic_vector(3 downto 0) := "1010";
  constant ANDOP: std_logic_vector(3 downto 0) := "1011";

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
      -- Inicializa os endereços:
tmp(0) := LDI&"00"&'0'&x"00";
tmp(1) := STA&"00"&'1'&x"20";
tmp(2) := STA&"00"&'1'&x"21";
tmp(3) := STA&"00"&'1'&x"22";
tmp(4) := STA&"00"&'1'&x"23";
tmp(5) := STA&"00"&'1'&x"24";
tmp(6) := STA&"00"&'1'&x"25";
tmp(7) := STA&"00"&'1'&x"00";
tmp(8) := STA&"00"&'1'&x"01";
tmp(9) := STA&"00"&'1'&x"02";
tmp(10) := STA&"00"&'0'&x"00";
tmp(11) := STA&"00"&'0'&x"01";
tmp(12) := STA&"00"&'0'&x"02";
tmp(13) := STA&"00"&'0'&x"03";
tmp(14) := STA&"00"&'0'&x"04";
tmp(15) := STA&"00"&'0'&x"05";
tmp(16) := STA&"00"&'0'&x"06";
tmp(17) := STA&"00"&'1'&x"ff";
tmp(18) := STA&"00"&'1'&x"fe";
tmp(19) := LDI&"00"&'0'&x"01";
tmp(20) := STA&"00"&'0'&x"0e";
tmp(22) := LDI&"00"&'0'&x"0a";
tmp(23) := STA&"00"&'0'&x"0f";
tmp(25) := LDI&"00"&'0'&x"00";
tmp(26) := STA&"00"&'0'&x"10";
tmp(28) := STA&"00"&'0'&x"08";
tmp(29) := STA&"00"&'0'&x"09";
tmp(30) := STA&"00"&'0'&x"0a";
tmp(31) := STA&"00"&'0'&x"0b";
tmp(32) := STA&"00"&'0'&x"0c";
tmp(33) := STA&"00"&'0'&x"0d";
tmp(38) := JSR&"00"&'0'&x"42";
tmp(40) := JSR&"00"&'1'&x"0e";
tmp(42) := LDA&"00"&'1'&x"60";
tmp(43) := ANDOP&"00"&'0'&x"0e";
tmp(44) := CEQ&"00"&'0'&x"06";
tmp(45) := JEQ&"00"&'0'&x"2f";
tmp(46) := JSR&"00"&'0'&x"57";
tmp(49) := LDA&"00"&'1'&x"61";
tmp(50) := ANDOP&"00"&'0'&x"0e";
tmp(51) := CEQ&"00"&'0'&x"06";
tmp(52) := JEQ&"00"&'0'&x"36";
tmp(53) := JSR&"00"&'0'&x"a9";
tmp(56) := LDA&"00"&'1'&x"64";
tmp(57) := ANDOP&"00"&'0'&x"0e";
tmp(58) := CEQ&"00"&'0'&x"06";
tmp(59) := JEQ&"00"&'0'&x"3d";
tmp(60) := JSR&"00"&'1'&x"39";
tmp(63) := JMP&"00"&'0'&x"24";
tmp(67) := LDA&"10"&'0'&x"00";
tmp(68) := STA&"10"&'1'&x"20";
tmp(69) := NOP&"00"&'0'&x"00";
tmp(70) := LDA&"10"&'0'&x"01";
tmp(71) := STA&"10"&'1'&x"21";
tmp(72) := NOP&"00"&'0'&x"00";
tmp(73) := LDA&"10"&'0'&x"02";
tmp(74) := STA&"10"&'1'&x"22";
tmp(75) := NOP&"00"&'0'&x"00";
tmp(76) := LDA&"10"&'0'&x"03";
tmp(77) := STA&"10"&'1'&x"23";
tmp(78) := NOP&"00"&'0'&x"00";
tmp(79) := LDA&"10"&'0'&x"04";
tmp(80) := STA&"10"&'1'&x"24";
tmp(81) := NOP&"00"&'0'&x"00";
tmp(82) := LDA&"10"&'0'&x"05";
tmp(83) := STA&"10"&'1'&x"25";
tmp(84) := RET&"00"&'0'&x"00";
tmp(88) := STA&"00"&'1'&x"ff";
tmp(89) := LDA&"00"&'0'&x"10";
tmp(90) := CEQ&"00"&'0'&x"0e";
tmp(91) := JEQ&"00"&'0'&x"a5";
tmp(93) := LDA&"00"&'0'&x"00";
tmp(94) := SOMA&"00"&'0'&x"0e";
tmp(95) := STA&"00"&'0'&x"00";
tmp(96) := CEQ&"00"&'0'&x"0f";
tmp(97) := JEQ&"00"&'0'&x"65";
tmp(98) := NOP&"00"&'0'&x"00";
tmp(99) := RET&"00"&'0'&x"00";
tmp(102) := LDI&"00"&'0'&x"00";
tmp(103) := STA&"00"&'0'&x"00";
tmp(104) := LDA&"00"&'0'&x"01";
tmp(105) := SOMA&"00"&'0'&x"0e";
tmp(106) := STA&"00"&'0'&x"01";
tmp(107) := CEQ&"00"&'0'&x"0f";
tmp(108) := JEQ&"00"&'0'&x"70";
tmp(109) := NOP&"00"&'0'&x"00";
tmp(110) := RET&"00"&'0'&x"00";
tmp(113) := LDI&"00"&'0'&x"00";
tmp(114) := STA&"00"&'0'&x"01";
tmp(115) := LDA&"00"&'0'&x"02";
tmp(116) := SOMA&"00"&'0'&x"0e";
tmp(117) := STA&"00"&'0'&x"02";
tmp(118) := CEQ&"00"&'0'&x"0f";
tmp(119) := JEQ&"00"&'0'&x"7b";
tmp(120) := NOP&"00"&'0'&x"00";
tmp(121) := RET&"00"&'0'&x"00";
tmp(124) := LDI&"00"&'0'&x"00";
tmp(125) := STA&"00"&'0'&x"02";
tmp(126) := LDA&"00"&'0'&x"03";
tmp(127) := SOMA&"00"&'0'&x"0e";
tmp(128) := STA&"00"&'0'&x"03";
tmp(129) := CEQ&"00"&'0'&x"0f";
tmp(130) := JEQ&"00"&'0'&x"86";
tmp(131) := NOP&"00"&'0'&x"00";
tmp(132) := RET&"00"&'0'&x"00";
tmp(135) := LDI&"00"&'0'&x"00";
tmp(136) := STA&"00"&'0'&x"03";
tmp(137) := LDA&"00"&'0'&x"04";
tmp(138) := SOMA&"00"&'0'&x"0e";
tmp(139) := STA&"00"&'0'&x"04";
tmp(140) := CEQ&"00"&'0'&x"0f";
tmp(141) := JEQ&"00"&'0'&x"91";
tmp(142) := NOP&"00"&'0'&x"00";
tmp(143) := RET&"00"&'0'&x"00";
tmp(146) := LDI&"00"&'0'&x"00";
tmp(147) := STA&"00"&'0'&x"04";
tmp(148) := LDA&"00"&'0'&x"05";
tmp(149) := SOMA&"00"&'0'&x"0e";
tmp(150) := STA&"00"&'0'&x"05";
tmp(151) := CEQ&"00"&'0'&x"0f";
tmp(152) := JEQ&"00"&'0'&x"9c";
tmp(153) := NOP&"00"&'0'&x"00";
tmp(154) := RET&"00"&'0'&x"00";
tmp(157) := LDI&"00"&'0'&x"00";
tmp(158) := STA&"00"&'0'&x"02";
tmp(160) := LDI&"00"&'0'&x"01";
tmp(161) := STA&"00"&'1'&x"02";
tmp(162) := STA&"00"&'0'&x"10";
tmp(166) := RET&"00"&'0'&x"00";
tmp(170) := STA&"00"&'1'&x"fe";
tmp(172) := LDI&"00"&'0'&x"01";
tmp(173) := STA&"00"&'1'&x"01";
tmp(174) := STA&"00"&'1'&x"02";
tmp(177) := LDI&"00"&'0'&x"01";
tmp(178) := STA&"00"&'1'&x"00";
tmp(179) := LDA&"00"&'1'&x"40";
tmp(180) := STA&"00"&'0'&x"08";
tmp(182) := LDA&"00"&'1'&x"61";
tmp(183) := ANDOP&"00"&'0'&x"0e";
tmp(184) := CEQ&"00"&'0'&x"06";
tmp(185) := JEQ&"00"&'0'&x"b0";
tmp(187) := LDI&"00"&'0'&x"00";
tmp(188) := STA&"00"&'1'&x"00";
tmp(189) := STA&"00"&'1'&x"fe";
tmp(192) := LDI&"00"&'0'&x"02";
tmp(193) := STA&"00"&'1'&x"00";
tmp(194) := LDA&"00"&'1'&x"40";
tmp(195) := STA&"00"&'0'&x"09";
tmp(197) := LDA&"00"&'1'&x"61";
tmp(198) := ANDOP&"00"&'0'&x"0e";
tmp(199) := CEQ&"00"&'0'&x"06";
tmp(200) := JEQ&"00"&'0'&x"bf";
tmp(202) := LDI&"00"&'0'&x"00";
tmp(203) := STA&"00"&'1'&x"00";
tmp(204) := STA&"00"&'1'&x"fe";
tmp(207) := LDI&"00"&'0'&x"04";
tmp(208) := STA&"00"&'1'&x"00";
tmp(209) := LDA&"00"&'1'&x"40";
tmp(210) := STA&"00"&'0'&x"0a";
tmp(212) := LDA&"00"&'1'&x"61";
tmp(213) := ANDOP&"00"&'0'&x"0e";
tmp(214) := CEQ&"00"&'0'&x"06";
tmp(215) := JEQ&"00"&'0'&x"ce";
tmp(217) := LDI&"00"&'0'&x"00";
tmp(218) := STA&"00"&'1'&x"00";
tmp(219) := STA&"00"&'1'&x"fe";
tmp(222) := LDI&"00"&'0'&x"08";
tmp(223) := STA&"00"&'1'&x"00";
tmp(224) := LDA&"00"&'1'&x"40";
tmp(225) := STA&"00"&'0'&x"0b";
tmp(227) := LDA&"00"&'1'&x"61";
tmp(228) := ANDOP&"00"&'0'&x"0e";
tmp(229) := CEQ&"00"&'0'&x"06";
tmp(230) := JEQ&"00"&'0'&x"dd";
tmp(232) := LDI&"00"&'0'&x"00";
tmp(233) := STA&"00"&'1'&x"00";
tmp(234) := STA&"00"&'1'&x"fe";
tmp(237) := LDI&"00"&'0'&x"10";
tmp(238) := STA&"00"&'1'&x"00";
tmp(239) := LDA&"00"&'1'&x"40";
tmp(240) := STA&"00"&'0'&x"0c";
tmp(242) := LDA&"00"&'1'&x"61";
tmp(243) := ANDOP&"00"&'0'&x"0e";
tmp(244) := CEQ&"00"&'0'&x"06";
tmp(245) := JEQ&"00"&'0'&x"ec";
tmp(247) := LDI&"00"&'0'&x"00";
tmp(248) := STA&"00"&'1'&x"00";
tmp(249) := STA&"00"&'1'&x"fe";
tmp(252) := LDI&"00"&'0'&x"20";
tmp(253) := STA&"00"&'1'&x"00";
tmp(254) := LDA&"00"&'1'&x"40";
tmp(255) := STA&"00"&'0'&x"0d";
tmp(257) := LDA&"00"&'1'&x"61";
tmp(258) := ANDOP&"00"&'0'&x"0e";
tmp(259) := CEQ&"00"&'0'&x"06";
tmp(260) := JEQ&"00"&'0'&x"fb";
tmp(262) := LDI&"00"&'0'&x"00";
tmp(263) := STA&"00"&'1'&x"00";
tmp(264) := STA&"00"&'1'&x"fe";
tmp(266) := STA&"00"&'1'&x"01";
tmp(267) := STA&"00"&'1'&x"02";
tmp(268) := JMP&"00"&'0'&x"24";
tmp(272) := LDA&"01"&'0'&x"05";
tmp(273) := CEQ&"01"&'0'&x"0d";
tmp(274) := JEQ&"00"&'1'&x"15";
tmp(275) := RET&"00"&'0'&x"00";
tmp(278) := LDA&"01"&'0'&x"04";
tmp(279) := CEQ&"01"&'0'&x"0c";
tmp(280) := JEQ&"00"&'1'&x"1b";
tmp(281) := RET&"00"&'0'&x"00";
tmp(284) := LDA&"01"&'0'&x"03";
tmp(285) := CEQ&"01"&'0'&x"0b";
tmp(286) := JEQ&"00"&'1'&x"21";
tmp(287) := RET&"00"&'0'&x"00";
tmp(290) := LDA&"01"&'0'&x"02";
tmp(291) := CEQ&"01"&'0'&x"0a";
tmp(292) := JEQ&"00"&'1'&x"27";
tmp(293) := RET&"00"&'0'&x"00";
tmp(296) := LDA&"01"&'0'&x"01";
tmp(297) := CEQ&"01"&'0'&x"09";
tmp(298) := JEQ&"00"&'1'&x"2d";
tmp(299) := RET&"00"&'0'&x"00";
tmp(302) := LDA&"01"&'0'&x"00";
tmp(303) := CEQ&"01"&'0'&x"08";
tmp(304) := JEQ&"00"&'1'&x"33";
tmp(305) := RET&"00"&'0'&x"00";
tmp(308) := LDI&"01"&'0'&x"01";
tmp(309) := STA&"01"&'0'&x"10";
tmp(310) := STA&"01"&'1'&x"01";
tmp(311) := RET&"00"&'0'&x"00";
tmp(314) := STA&"00"&'1'&x"fc";
tmp(315) := LDI&"00"&'0'&x"00";
tmp(316) := STA&"00"&'0'&x"00";
tmp(317) := STA&"00"&'0'&x"01";
tmp(318) := STA&"00"&'0'&x"02";
tmp(319) := STA&"00"&'0'&x"03";
tmp(320) := STA&"00"&'0'&x"04";
tmp(321) := STA&"00"&'0'&x"05";
tmp(322) := STA&"00"&'0'&x"10";
tmp(323) := STA&"00"&'1'&x"01";
tmp(324) := STA&"00"&'1'&x"02";
tmp(325) := STA&"00"&'1'&x"00";
tmp(327) := RET&"00"&'0'&x"00";





        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;